package ahb_apb_pkg;

    import uvm_pkg::*;
	
        `include "uvm_macros.svh"
	`include "ahb_xtns.sv"
	`include "ahb_agt_config.sv"
	`include "apb_agt_config.sv"
	`include "ahb_apb_env_config.sv"

	`include "ahb_driver.sv"
	`include "ahb_monitor.sv"
	`include "ahb_sequencer.sv"
	`include "ahb_agt.sv"
	`include "ahb_agt_top.sv"
	`include "ahb_seq.sv"

	`include "apb_xtns.sv"
  `include "apb_driver.sv"
	`include "apb_monitor.sv"
	`include "apb_sequencer.sv"
	`include "apb_agt.sv"
	`include "apb_agt_top.sv"
	`include "apb_seq.sv"
	
  
  `include "ahb_apb_v_sequencer.sv"
  `include "ahb_apb_v_sequence.sv"
  `include "ahb_apb_scoreboard.sv"
	`include "ahb_apb_env.sv"
	`include "ahb_apb_test.sv"
	
endpackage
